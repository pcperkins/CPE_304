-- Contact me if you want the code.
